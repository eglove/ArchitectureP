library verilog;
use verilog.vl_types.all;
entity top_tb is
    generic(
        CLK_CYCLE       : integer := 50
    );
end top_tb;

library verilog;
use verilog.vl_types.all;
entity \32-bitProcessor\ is
end \32-bitProcessor\;

`timescale 1ns/1ps

module signext#(parameter IN=5, OUT=10)
(
	input [IN-1:0] din,
	output [OUT-1:0] dout
);

endmodule
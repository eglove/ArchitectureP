module controller (input clk,reset,
               input [5:0] op, funct,
				   output memtoreg, memwrite,
				   output alusrca,
				   output [1:0] alusrcb,
				   output regdst, regwrite,
				   output jump,signext,
				   output [3:0] alucontrol,
					output branch,
					output PCWriteCond,PCWrite,
					output IorD,IRWrite,
					output [1:0] pcsrc
); //controller signals

	wire [2:0] aluop;        //determine what the alu is to do
	wire [15:0] state;         //FSM
	maindec md (clk,reset,op, memtoreg, memwrite, branch,
	alusrca,alusrcb, regdst, regwrite, jump,signext,
	aluop,PCWriteCond,PCWrite,IorD,IRWrite,state,pcsrc);       //main decoder produces main signales
	//alu decoder produces the direct signal to control alu
	aludec ad (funct, aluop, alucontrol);      
endmodule
